`timescale 1ns/10ps
module Control_tb();

	reg [31:0] in;
	wire [22:0] out;

	Control DUT(
		.in(in),
		.out(out)
	);

	initial begin
		in = 32'b0;
		
		#10 in = 32'b000101_00000_00001_0011_0000_0000_0000; //LW
		#10 in = 32'b000110_00000_00001_0000_0000_0000_0000; //SW
		#10 in = 32'b000100_00000_00001_00010_01010_100000;  //ADD
		#10 in = 32'b000100_00000_00001_00010_01010_100010;  //SUB
		#10 in = 32'b000100_00000_00001_00010_01010_110010;  //MUL
		#10 in = 32'b000100_00000_00001_00010_01010_100100;  //AND
		#10 in = 32'b000100_00000_00001_00010_01010_100101;  //OR
	
	//	#10 in = 32'b001111_00000_00010_0001_0100_0000_0000; //LW
	//#10 in = 32'b010000_00000_01101_0001_1000_0000_0000; //SW
	//	#10 in = 32'b000100_00101_00111_01011_01010_100000;   //ADD
	//	#10 in = 32'b000100_01100_01011_01101_01010_100010;  //SUB
	//	#10 in = 32'b000100_00010_00011_01100_01010_110010;  //MUL
	//	#10 in = 32'b001110_00000_00001_00010_01010_100100;  //AND
	//	#10 in = 32'b001110_00000_00001_00010_01010_100101;  //OR
		#10 $stop;
		
	end
	
endmodule 